`timescale 1ns / 1ps

module MUX2s32b(
    );


endmodule
