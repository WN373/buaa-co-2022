module EX2MEM (
    
);

endmodule