module hazard(
    input [31:0] D_ins, E_ins, M_ins,

);

endmodule