module Controller(
    input [5:0] optCode, funcCode
    output reg_write_enable, mem_write_enable, 
    output [3:0] alu_op, ext_op,
    output [2:0] nPC_sel
);
    

endmodule